library verilog;
use verilog.vl_types.all;
entity tb_aluCtrl is
end tb_aluCtrl;
