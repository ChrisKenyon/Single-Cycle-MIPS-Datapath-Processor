library verilog;
use verilog.vl_types.all;
entity tb_ctrlUnit is
end tb_ctrlUnit;
